module not1(s,y);
input s;
output y;
assign y = ~s;
endmodule
